    Mac OS X            	   2   �      �                                      ATTR       �   �   *                  �     com.apple.lastuseddate#PS       �     com.dropbox.attrs    �WO`    wZ/    

`,���f�       ����