    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

�5 ���b�       ����