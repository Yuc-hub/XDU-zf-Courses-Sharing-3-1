    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

ԇ�hr
�p       ���