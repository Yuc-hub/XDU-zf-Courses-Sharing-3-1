    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

8�rj߿l�       ����