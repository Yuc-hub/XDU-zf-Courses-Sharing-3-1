LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


entity ADDC4 is 
port (
			I1, I2: in std_logic_vector(3 downto 0);
			CIN : in std_logic;
			SUM  : out std_logic_vector(3 downto 0); 
			COUT : out  std_logic );
end entity ADDC4;



architecture STRUCT of ADDC4 is
begin
	
	 
end architecture STRUCT;
