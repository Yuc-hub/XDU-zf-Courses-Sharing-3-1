    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

|�?(橧        �ѡ�