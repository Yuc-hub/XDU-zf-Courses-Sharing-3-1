-- Squelette pour l'exercice carte m�moire

library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.numeric_std.all;

entity Board is
  generic (ChipAddressSize : integer);
  port (Address: in Std_logic_vector(7 downto 0);
        Data: inout Std_logic_vector(15 downto 0);
        nWE, nOE: in Std_logic);
end entity Board;

architecture Struct of Board is
   signal A : Std_logic_vector(Address'high-ChipAddressSize downto 0);
   signal B : Std_logic_vector(ChipAddressSize-1 downto 0);
   signal C : Std_logic_vector(2**(Address'high-ChipAddressSize+1)-1 downto 0);
begin
   A <= Address(Address'high downto ChipAddressSize);
   B <= Address(ChipAddressSize-1 downto 0);
C <= (others => '0');
C(to_integer(unsigned(A))) <= '1';

L1: for I in 0 to 2**(Address'high-ChipAddressSize+1)-1 generate
	U1 : entity work.ramchip generic map(4, 16)
        port map(nCS => C(I), Address => B, nWE => nWE, nOE => nOE, Data => Data);
end generate;
end architecture Struct;