-- Squelette pour l'exercice sur les machines � �tats

library IEEE;
use IEEE.STD_LOGIC_1164.all;                             
                                                         
entity FSM is                                            
								  port (	Clk :	in 	STD_LOGIC;                          
								  			nRst: in 	STD_LOGIC;                          
								       	Start_Stop, Clear:	in 	STD_LOGIC;           
								        	Cnt_En, Cnt_Rst: 		out 	STD_LOGIC);          
end entity;                                              
                                                         
architecture RTL of FSm is                               
begin                                                    
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
                                                         
end architecture;
