    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

1X��W\     �͉��